magic
tech scmos
timestamp 1695044485
<< nwell >>
rect -7 -5 9 6
<< polysilicon >>
rect -1 4 1 6
rect -1 -9 1 -3
rect -4 -12 1 -9
rect -1 -17 1 -12
rect -1 -26 1 -23
<< ndiffusion >>
rect -7 -18 -1 -17
rect -7 -23 -6 -18
rect -2 -23 -1 -18
rect 1 -18 5 -17
rect 1 -23 2 -18
<< pdiffusion >>
rect -6 1 -1 4
rect -2 -3 -1 1
rect 1 1 6 4
rect 1 -3 2 1
<< metal1 >>
rect -6 17 5 19
rect -2 13 5 17
rect -6 8 5 13
rect -6 1 -2 8
rect 2 1 5 3
rect 2 -8 5 -3
rect 2 -12 8 -8
rect 2 -18 5 -12
rect -6 -29 -2 -23
rect -6 -32 5 -29
rect -2 -36 5 -32
<< ntransistor >>
rect -1 -23 1 -17
<< ptransistor >>
rect -1 -3 1 4
<< ndcontact >>
rect -6 -23 -2 -18
rect 2 -23 6 -18
<< pdcontact >>
rect -6 -3 -2 1
rect 2 -3 6 1
<< psubstratepcontact >>
rect -6 13 -2 17
<< nsubstratencontact >>
rect -6 -36 -2 -32
<< labels >>
rlabel metal1 2 -12 8 -8 7 out
rlabel polysilicon -4 -12 -1 -9 3 in
rlabel metal1 -1 8 3 11 5 vdd
rlabel metal1 -1 -32 3 -29 1 gnd
<< end >>
